--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   12:46:58 02/15/2016
-- Design Name:   
-- Module Name:   U:/Project-1-Datapath-Design-Part-A-2/mux8_16bit_tb.vhd
-- Project Name:  Project-1-Datapath-Design-Part-A-2
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: mux8_16bit
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY mux8_16bit_tb IS
END mux8_16bit_tb;
 
ARCHITECTURE behavior OF mux8_16bit_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT mux8_16bit
    PORT(
         in0 : IN  std_logic_vector(15 downto 0);
         in1 : IN  std_logic_vector(15 downto 0);
         in2 : IN  std_logic_vector(15 downto 0);
         in3 : IN  std_logic_vector(15 downto 0);
         in4 : IN  std_logic_vector(15 downto 0);
         in5 : IN  std_logic_vector(15 downto 0);
         in6 : IN  std_logic_vector(15 downto 0);
         in7 : IN  std_logic_vector(15 downto 0);
         s0 : IN  std_logic;
         s1 : IN  std_logic;
         s2 : IN  std_logic;
         z : OUT  std_logic_vector(15 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal in0 : std_logic_vector(15 downto 0) := (others => '0');
   signal in1 : std_logic_vector(15 downto 0) := (others => '0');
   signal in2 : std_logic_vector(15 downto 0) := (others => '0');
   signal in3 : std_logic_vector(15 downto 0) := (others => '0');
   signal in4 : std_logic_vector(15 downto 0) := (others => '0');
   signal in5 : std_logic_vector(15 downto 0) := (others => '0');
   signal in6 : std_logic_vector(15 downto 0) := (others => '0');
   signal in7 : std_logic_vector(15 downto 0) := (others => '0');
   signal s0 : std_logic := '0';
   signal s1 : std_logic := '0';
   signal s2 : std_logic := '0';

 	--Outputs
   signal z : std_logic_vector(15 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: mux8_16bit PORT MAP (
          in0 => in0,
          in1 => in1,
          in2 => in2,
          in3 => in3,
          in4 => in4,
          in5 => in5,
          in6 => in6,
          in7 => in7,
          s0 => s0,
          s1 => s1,
          s2 => s2,
          z => z
        );

   -- Stimulus process
   stim_proc: process
   begin		
	
		in0 <=	X"df23";
		in1 <=	X"f87d";
		in2 <=	X"ffff";
		in3 <=	X"90ac";
		in4 <=	X"7ef6";
		in5 <=	X"f91a";
		in6 <=	X"3cd4";
		in7 <=	X"b4a2";
		
		s0 <= '0';
		s1 <= '0';
		s2 <= '0';
	
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      s0 <= '0';
		s1 <= '0';
		s2 <= '1';
		
		wait for 100 ns;
		
		s0 <= '0';
		s1 <= '1';
		s2 <= '0';
		
		wait for 100 ns;
		
		s0 <= '0';
		s1 <= '1';
		s2 <= '1';
		
		wait for 100 ns;
		
		s0 <= '1';
		s1 <= '0';
		s2 <= '0';
		
		wait for 100 ns;
		
		s0 <= '1';
		s1 <= '0';
		s2 <= '1';
		
		wait for 100 ns;
		
		s0 <= '1';
		s1 <= '1';
		s2 <= '0';
		
		wait for 100 ns;
		
		s0 <= '1';
		s1 <= '1';
		s2 <= '1';

      wait;
   end process;

END;
